`default_nettype none

module execute_stage(
    input wire i_clk, i_reset,
);



endmodule : execute