`default_nettype none

module execute(
    input wire i_clk, i_reset,
);



endmodule : execute